module ICache();

endmodule