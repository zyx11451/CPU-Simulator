module register (
    
);

  reg [31:0] reg_value[31:0];
  
endmodule  //register

